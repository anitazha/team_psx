`define SCREEN_H 9'd480
`define SCREEN_W 10'd640
